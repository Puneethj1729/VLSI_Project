magic
tech scmos
timestamp 1608657425
<< pwell >>
rect -110 239 -84 262
rect -111 135 -85 158
rect 8 139 69 171
rect 148 139 209 171
rect 288 139 349 171
rect 435 139 496 171
rect 569 139 630 171
rect 706 139 767 171
rect 845 139 906 171
rect 980 139 1041 171
rect -109 26 -83 49
<< nwell >>
rect -110 278 -84 319
rect -111 174 -85 215
rect 8 208 69 237
rect 148 208 209 237
rect 288 208 349 237
rect 435 208 496 237
rect 569 208 630 237
rect 706 208 767 237
rect 845 208 906 237
rect 980 208 1041 237
rect -109 65 -83 106
<< polysilicon >>
rect -98 309 -96 311
rect -98 261 -96 279
rect -98 247 -96 249
rect 18 224 20 226
rect 28 224 30 226
rect 37 224 39 226
rect 57 225 59 227
rect -99 205 -97 207
rect -99 157 -97 175
rect 18 170 20 209
rect 28 170 30 209
rect 37 170 39 209
rect 158 224 160 226
rect 168 224 170 226
rect 177 224 179 226
rect 197 225 199 227
rect 57 162 59 208
rect 158 170 160 209
rect 168 170 170 209
rect 177 170 179 209
rect 298 224 300 226
rect 308 224 310 226
rect 317 224 319 226
rect 337 225 339 227
rect 57 154 59 156
rect 197 162 199 208
rect 298 170 300 209
rect 308 170 310 209
rect 317 170 319 209
rect 445 224 447 226
rect 455 224 457 226
rect 464 224 466 226
rect 484 225 486 227
rect 197 154 199 156
rect 337 162 339 208
rect 445 170 447 209
rect 455 170 457 209
rect 464 170 466 209
rect 579 224 581 226
rect 589 224 591 226
rect 598 224 600 226
rect 618 225 620 227
rect 337 154 339 156
rect 484 162 486 208
rect 579 170 581 209
rect 589 170 591 209
rect 598 170 600 209
rect 716 224 718 226
rect 726 224 728 226
rect 735 224 737 226
rect 755 225 757 227
rect 484 154 486 156
rect 618 162 620 208
rect 716 170 718 209
rect 726 170 728 209
rect 735 170 737 209
rect 855 224 857 226
rect 865 224 867 226
rect 874 224 876 226
rect 894 225 896 227
rect 618 154 620 156
rect 755 162 757 208
rect 855 170 857 209
rect 865 170 867 209
rect 874 170 876 209
rect 990 224 992 226
rect 1000 224 1002 226
rect 1009 224 1011 226
rect 1029 225 1031 227
rect 755 154 757 156
rect 894 162 896 208
rect 990 170 992 209
rect 1000 170 1002 209
rect 1009 170 1011 209
rect 894 154 896 156
rect 1029 162 1031 208
rect 1029 154 1031 156
rect 18 150 20 152
rect 28 150 30 152
rect 37 150 39 152
rect 158 150 160 152
rect 168 150 170 152
rect 177 150 179 152
rect 298 150 300 152
rect 308 150 310 152
rect 317 150 319 152
rect 445 150 447 152
rect 455 150 457 152
rect 464 150 466 152
rect 579 150 581 152
rect 589 150 591 152
rect 598 150 600 152
rect 716 150 718 152
rect 726 150 728 152
rect 735 150 737 152
rect 855 150 857 152
rect 865 150 867 152
rect 874 150 876 152
rect 990 150 992 152
rect 1000 150 1002 152
rect 1009 150 1011 152
rect -99 143 -97 145
rect -97 96 -95 98
rect -97 48 -95 66
rect -97 34 -95 36
<< ndiffusion >>
rect -99 257 -98 261
rect -103 253 -98 257
rect -99 249 -98 253
rect -96 257 -95 261
rect -96 253 -91 257
rect -96 249 -95 253
rect 17 166 18 170
rect 13 163 18 166
rect 17 159 18 163
rect -100 153 -99 157
rect -104 149 -99 153
rect -100 145 -99 149
rect -97 153 -96 157
rect -97 149 -92 153
rect 13 156 18 159
rect 17 152 18 156
rect 20 152 28 170
rect 30 152 37 170
rect 39 166 40 170
rect 39 163 44 166
rect 39 159 40 163
rect 157 166 158 170
rect 153 163 158 166
rect 39 156 44 159
rect 52 161 57 162
rect 56 157 57 161
rect 52 156 57 157
rect 59 161 64 162
rect 59 157 60 161
rect 59 156 64 157
rect 157 159 158 163
rect 153 156 158 159
rect 39 152 40 156
rect 157 152 158 156
rect 160 152 168 170
rect 170 152 177 170
rect 179 166 180 170
rect 179 163 184 166
rect 179 159 180 163
rect 297 166 298 170
rect 293 163 298 166
rect 179 156 184 159
rect 192 161 197 162
rect 196 157 197 161
rect 192 156 197 157
rect 199 161 204 162
rect 199 157 200 161
rect 199 156 204 157
rect 297 159 298 163
rect 293 156 298 159
rect 179 152 180 156
rect 297 152 298 156
rect 300 152 308 170
rect 310 152 317 170
rect 319 166 320 170
rect 319 163 324 166
rect 319 159 320 163
rect 444 166 445 170
rect 440 163 445 166
rect 319 156 324 159
rect 332 161 337 162
rect 336 157 337 161
rect 332 156 337 157
rect 339 161 344 162
rect 339 157 340 161
rect 339 156 344 157
rect 444 159 445 163
rect 440 156 445 159
rect 319 152 320 156
rect 444 152 445 156
rect 447 152 455 170
rect 457 152 464 170
rect 466 166 467 170
rect 466 163 471 166
rect 466 159 467 163
rect 578 166 579 170
rect 574 163 579 166
rect 466 156 471 159
rect 479 161 484 162
rect 483 157 484 161
rect 479 156 484 157
rect 486 161 491 162
rect 486 157 487 161
rect 486 156 491 157
rect 578 159 579 163
rect 574 156 579 159
rect 466 152 467 156
rect 578 152 579 156
rect 581 152 589 170
rect 591 152 598 170
rect 600 166 601 170
rect 600 163 605 166
rect 600 159 601 163
rect 715 166 716 170
rect 711 163 716 166
rect 600 156 605 159
rect 613 161 618 162
rect 617 157 618 161
rect 613 156 618 157
rect 620 161 625 162
rect 620 157 621 161
rect 620 156 625 157
rect 715 159 716 163
rect 711 156 716 159
rect 600 152 601 156
rect 715 152 716 156
rect 718 152 726 170
rect 728 152 735 170
rect 737 166 738 170
rect 737 163 742 166
rect 737 159 738 163
rect 854 166 855 170
rect 850 163 855 166
rect 737 156 742 159
rect 750 161 755 162
rect 754 157 755 161
rect 750 156 755 157
rect 757 161 762 162
rect 757 157 758 161
rect 757 156 762 157
rect 854 159 855 163
rect 850 156 855 159
rect 737 152 738 156
rect 854 152 855 156
rect 857 152 865 170
rect 867 152 874 170
rect 876 166 877 170
rect 876 163 881 166
rect 876 159 877 163
rect 989 166 990 170
rect 985 163 990 166
rect 876 156 881 159
rect 889 161 894 162
rect 893 157 894 161
rect 889 156 894 157
rect 896 161 901 162
rect 896 157 897 161
rect 896 156 901 157
rect 989 159 990 163
rect 985 156 990 159
rect 876 152 877 156
rect 989 152 990 156
rect 992 152 1000 170
rect 1002 152 1009 170
rect 1011 166 1012 170
rect 1011 163 1016 166
rect 1011 159 1012 163
rect 1011 156 1016 159
rect 1024 161 1029 162
rect 1028 157 1029 161
rect 1024 156 1029 157
rect 1031 161 1036 162
rect 1031 157 1032 161
rect 1031 156 1036 157
rect 1011 152 1012 156
rect -97 145 -96 149
rect -98 44 -97 48
rect -102 40 -97 44
rect -98 36 -97 40
rect -95 44 -94 48
rect -95 40 -90 44
rect -95 36 -94 40
<< pdiffusion >>
rect -103 308 -98 309
rect -99 304 -98 308
rect -103 299 -98 304
rect -99 295 -98 299
rect -103 291 -98 295
rect -99 287 -98 291
rect -103 283 -98 287
rect -99 279 -98 283
rect -96 308 -91 309
rect -96 304 -95 308
rect -96 299 -91 304
rect -96 295 -95 299
rect -96 291 -91 295
rect -96 287 -95 291
rect -96 283 -91 287
rect -96 279 -95 283
rect 52 224 57 225
rect 17 220 18 224
rect 13 213 18 220
rect 17 209 18 213
rect 20 220 22 224
rect 26 220 28 224
rect 20 213 28 220
rect 20 209 22 213
rect 26 209 28 213
rect 30 220 32 224
rect 36 220 37 224
rect 30 213 37 220
rect 30 209 32 213
rect 36 209 37 213
rect 39 220 40 224
rect 39 213 44 220
rect 39 209 40 213
rect 56 220 57 224
rect 52 218 57 220
rect 56 214 57 218
rect 52 212 57 214
rect -104 204 -99 205
rect -100 200 -99 204
rect -104 195 -99 200
rect -100 191 -99 195
rect -104 187 -99 191
rect -100 183 -99 187
rect -104 179 -99 183
rect -100 175 -99 179
rect -97 204 -92 205
rect -97 200 -96 204
rect -97 195 -92 200
rect -97 191 -96 195
rect -97 187 -92 191
rect -97 183 -96 187
rect -97 179 -92 183
rect -97 175 -96 179
rect 56 208 57 212
rect 59 224 64 225
rect 192 224 197 225
rect 59 220 60 224
rect 59 218 64 220
rect 59 214 60 218
rect 59 212 64 214
rect 59 208 60 212
rect 157 220 158 224
rect 153 213 158 220
rect 157 209 158 213
rect 160 220 162 224
rect 166 220 168 224
rect 160 213 168 220
rect 160 209 162 213
rect 166 209 168 213
rect 170 220 172 224
rect 176 220 177 224
rect 170 213 177 220
rect 170 209 172 213
rect 176 209 177 213
rect 179 220 180 224
rect 179 213 184 220
rect 179 209 180 213
rect 196 220 197 224
rect 192 218 197 220
rect 196 214 197 218
rect 192 212 197 214
rect 196 208 197 212
rect 199 224 204 225
rect 332 224 337 225
rect 199 220 200 224
rect 199 218 204 220
rect 199 214 200 218
rect 199 212 204 214
rect 199 208 200 212
rect 297 220 298 224
rect 293 213 298 220
rect 297 209 298 213
rect 300 220 302 224
rect 306 220 308 224
rect 300 213 308 220
rect 300 209 302 213
rect 306 209 308 213
rect 310 220 312 224
rect 316 220 317 224
rect 310 213 317 220
rect 310 209 312 213
rect 316 209 317 213
rect 319 220 320 224
rect 319 213 324 220
rect 319 209 320 213
rect 336 220 337 224
rect 332 218 337 220
rect 336 214 337 218
rect 332 212 337 214
rect 336 208 337 212
rect 339 224 344 225
rect 479 224 484 225
rect 339 220 340 224
rect 339 218 344 220
rect 339 214 340 218
rect 339 212 344 214
rect 339 208 340 212
rect 444 220 445 224
rect 440 213 445 220
rect 444 209 445 213
rect 447 220 449 224
rect 453 220 455 224
rect 447 213 455 220
rect 447 209 449 213
rect 453 209 455 213
rect 457 220 459 224
rect 463 220 464 224
rect 457 213 464 220
rect 457 209 459 213
rect 463 209 464 213
rect 466 220 467 224
rect 466 213 471 220
rect 466 209 467 213
rect 483 220 484 224
rect 479 218 484 220
rect 483 214 484 218
rect 479 212 484 214
rect 483 208 484 212
rect 486 224 491 225
rect 613 224 618 225
rect 486 220 487 224
rect 486 218 491 220
rect 486 214 487 218
rect 486 212 491 214
rect 486 208 487 212
rect 578 220 579 224
rect 574 213 579 220
rect 578 209 579 213
rect 581 220 583 224
rect 587 220 589 224
rect 581 213 589 220
rect 581 209 583 213
rect 587 209 589 213
rect 591 220 593 224
rect 597 220 598 224
rect 591 213 598 220
rect 591 209 593 213
rect 597 209 598 213
rect 600 220 601 224
rect 600 213 605 220
rect 600 209 601 213
rect 617 220 618 224
rect 613 218 618 220
rect 617 214 618 218
rect 613 212 618 214
rect 617 208 618 212
rect 620 224 625 225
rect 750 224 755 225
rect 620 220 621 224
rect 620 218 625 220
rect 620 214 621 218
rect 620 212 625 214
rect 620 208 621 212
rect 715 220 716 224
rect 711 213 716 220
rect 715 209 716 213
rect 718 220 720 224
rect 724 220 726 224
rect 718 213 726 220
rect 718 209 720 213
rect 724 209 726 213
rect 728 220 730 224
rect 734 220 735 224
rect 728 213 735 220
rect 728 209 730 213
rect 734 209 735 213
rect 737 220 738 224
rect 737 213 742 220
rect 737 209 738 213
rect 754 220 755 224
rect 750 218 755 220
rect 754 214 755 218
rect 750 212 755 214
rect 754 208 755 212
rect 757 224 762 225
rect 889 224 894 225
rect 757 220 758 224
rect 757 218 762 220
rect 757 214 758 218
rect 757 212 762 214
rect 757 208 758 212
rect 854 220 855 224
rect 850 213 855 220
rect 854 209 855 213
rect 857 220 859 224
rect 863 220 865 224
rect 857 213 865 220
rect 857 209 859 213
rect 863 209 865 213
rect 867 220 869 224
rect 873 220 874 224
rect 867 213 874 220
rect 867 209 869 213
rect 873 209 874 213
rect 876 220 877 224
rect 876 213 881 220
rect 876 209 877 213
rect 893 220 894 224
rect 889 218 894 220
rect 893 214 894 218
rect 889 212 894 214
rect 893 208 894 212
rect 896 224 901 225
rect 1024 224 1029 225
rect 896 220 897 224
rect 896 218 901 220
rect 896 214 897 218
rect 896 212 901 214
rect 896 208 897 212
rect 989 220 990 224
rect 985 213 990 220
rect 989 209 990 213
rect 992 220 994 224
rect 998 220 1000 224
rect 992 213 1000 220
rect 992 209 994 213
rect 998 209 1000 213
rect 1002 220 1004 224
rect 1008 220 1009 224
rect 1002 213 1009 220
rect 1002 209 1004 213
rect 1008 209 1009 213
rect 1011 220 1012 224
rect 1011 213 1016 220
rect 1011 209 1012 213
rect 1028 220 1029 224
rect 1024 218 1029 220
rect 1028 214 1029 218
rect 1024 212 1029 214
rect 1028 208 1029 212
rect 1031 224 1036 225
rect 1031 220 1032 224
rect 1031 218 1036 220
rect 1031 214 1032 218
rect 1031 212 1036 214
rect 1031 208 1032 212
rect -102 95 -97 96
rect -98 91 -97 95
rect -102 86 -97 91
rect -98 82 -97 86
rect -102 78 -97 82
rect -98 74 -97 78
rect -102 70 -97 74
rect -98 66 -97 70
rect -95 95 -90 96
rect -95 91 -94 95
rect -95 86 -90 91
rect -95 82 -94 86
rect -95 78 -90 82
rect -95 74 -94 78
rect -95 70 -90 74
rect -95 66 -94 70
<< metal1 >>
rect -106 314 -99 318
rect -95 314 -88 318
rect -84 314 -60 318
rect -103 308 -99 314
rect -103 299 -99 304
rect -103 291 -99 295
rect -103 283 -99 287
rect -95 308 -91 309
rect -95 299 -91 304
rect -95 291 -91 295
rect -95 283 -91 287
rect -95 272 -91 279
rect -56 292 129 296
rect 133 292 273 296
rect 277 292 410 296
rect -56 272 -52 292
rect -155 268 -102 272
rect -95 268 -52 272
rect -155 -8 -151 268
rect -95 261 -91 268
rect -103 253 -99 257
rect -95 253 -91 257
rect -103 244 -99 249
rect -126 240 -110 244
rect -106 240 -99 244
rect -95 240 -88 244
rect -107 210 -100 214
rect -96 210 -89 214
rect -85 210 -60 214
rect -104 204 -100 210
rect -104 195 -100 200
rect -104 187 -100 191
rect -104 179 -100 183
rect -96 204 -92 205
rect -96 195 -92 200
rect -12 198 -8 292
rect 8 276 108 280
rect 112 276 554 280
rect 558 276 685 280
rect 8 260 263 264
rect 267 260 543 264
rect 547 260 798 264
rect 12 230 16 234
rect 20 230 24 234
rect 28 230 32 234
rect 36 230 40 234
rect 44 230 48 234
rect 22 224 26 230
rect 40 224 44 230
rect 13 213 17 220
rect 22 213 26 220
rect 32 213 36 220
rect 40 213 44 220
rect 52 224 56 234
rect 60 230 64 234
rect 68 230 76 234
rect 80 230 148 234
rect 152 230 156 234
rect 160 230 164 234
rect 168 230 172 234
rect 176 230 180 234
rect 184 230 188 234
rect 52 218 56 220
rect 52 212 56 214
rect 13 206 17 209
rect 32 206 36 209
rect 60 224 64 225
rect 162 224 166 230
rect 180 224 184 230
rect 60 218 64 220
rect 60 212 64 214
rect 13 202 47 206
rect -12 194 14 198
rect 43 191 47 202
rect 60 191 64 208
rect 153 213 157 220
rect 162 213 166 220
rect 172 213 176 220
rect 180 213 184 220
rect 192 224 196 234
rect 200 230 204 234
rect 208 230 288 234
rect 292 230 296 234
rect 300 230 304 234
rect 308 230 312 234
rect 316 230 320 234
rect 324 230 328 234
rect 192 218 196 220
rect 192 212 196 214
rect 153 206 157 209
rect 172 206 176 209
rect 200 224 204 225
rect 302 224 306 230
rect 320 224 324 230
rect 200 218 204 220
rect 200 212 204 214
rect 153 202 187 206
rect 133 194 154 198
rect 183 191 187 202
rect 200 191 204 208
rect 293 213 297 220
rect 302 213 306 220
rect 312 213 316 220
rect 320 213 324 220
rect 332 224 336 234
rect 340 230 344 234
rect 348 230 435 234
rect 439 230 443 234
rect 447 230 451 234
rect 455 230 459 234
rect 463 230 467 234
rect 471 230 475 234
rect 332 218 336 220
rect 332 212 336 214
rect 293 206 297 209
rect 312 206 316 209
rect 340 224 344 225
rect 449 224 453 230
rect 467 224 471 230
rect 340 218 344 220
rect 340 212 344 214
rect 293 202 327 206
rect 277 194 294 198
rect 323 191 327 202
rect 340 191 344 208
rect 440 213 444 220
rect 449 213 453 220
rect 459 213 463 220
rect 467 213 471 220
rect 479 224 483 234
rect 487 230 491 234
rect 495 230 569 234
rect 573 230 577 234
rect 581 230 585 234
rect 589 230 593 234
rect 597 230 601 234
rect 605 230 609 234
rect 479 218 483 220
rect 479 212 483 214
rect 440 206 444 209
rect 459 206 463 209
rect 487 224 491 225
rect 583 224 587 230
rect 601 224 605 230
rect 487 218 491 220
rect 487 212 491 214
rect 440 202 474 206
rect 414 194 441 198
rect 470 191 474 202
rect 487 191 491 208
rect 574 213 578 220
rect 583 213 587 220
rect 593 213 597 220
rect 601 213 605 220
rect 613 224 617 234
rect 621 230 625 234
rect 629 230 706 234
rect 710 230 714 234
rect 718 230 722 234
rect 726 230 730 234
rect 734 230 738 234
rect 742 230 746 234
rect 613 218 617 220
rect 613 212 617 214
rect 574 206 578 209
rect 593 206 597 209
rect 621 224 625 225
rect 720 224 724 230
rect 738 224 742 230
rect 621 218 625 220
rect 621 212 625 214
rect 574 202 608 206
rect 535 194 575 198
rect 604 191 608 202
rect 621 191 625 208
rect 711 213 715 220
rect 720 213 724 220
rect 730 213 734 220
rect 738 213 742 220
rect 750 224 754 234
rect 758 230 762 234
rect 766 230 845 234
rect 849 230 853 234
rect 857 230 861 234
rect 865 230 869 234
rect 873 230 877 234
rect 881 230 885 234
rect 750 218 754 220
rect 750 212 754 214
rect 711 206 715 209
rect 730 206 734 209
rect 758 224 762 225
rect 859 224 863 230
rect 877 224 881 230
rect 758 218 762 220
rect 758 212 762 214
rect 711 202 745 206
rect 673 194 712 198
rect 741 191 745 202
rect 758 191 762 208
rect 850 213 854 220
rect 859 213 863 220
rect 869 213 873 220
rect 877 213 881 220
rect 889 224 893 234
rect 897 230 901 234
rect 905 230 980 234
rect 984 230 988 234
rect 992 230 996 234
rect 1000 230 1004 234
rect 1008 230 1012 234
rect 1016 230 1020 234
rect 889 218 893 220
rect 889 212 893 214
rect 850 206 854 209
rect 869 206 873 209
rect 897 224 901 225
rect 994 224 998 230
rect 1012 224 1016 230
rect 897 218 901 220
rect 897 212 901 214
rect 850 202 884 206
rect 819 194 851 198
rect 880 191 884 202
rect 897 191 901 208
rect 985 213 989 220
rect 994 213 998 220
rect 1004 213 1008 220
rect 1012 213 1016 220
rect 1024 224 1028 234
rect 1032 230 1036 234
rect 1040 230 1041 234
rect 1024 218 1028 220
rect 1024 212 1028 214
rect 985 206 989 209
rect 1004 206 1008 209
rect 1032 224 1036 225
rect 1032 218 1036 220
rect 1032 212 1036 214
rect 985 202 1019 206
rect 974 194 986 198
rect 1015 191 1019 202
rect 1032 191 1036 208
rect -96 187 -92 191
rect -96 179 -92 183
rect -96 168 -92 175
rect -27 187 24 191
rect 43 187 53 191
rect 60 187 69 191
rect 112 187 164 191
rect 183 187 193 191
rect 200 187 209 191
rect 254 187 304 191
rect 323 187 333 191
rect 340 187 349 191
rect 402 187 451 191
rect 470 187 480 191
rect 487 187 496 191
rect 558 187 585 191
rect 604 187 614 191
rect 621 187 630 191
rect 689 187 722 191
rect 741 187 751 191
rect 758 187 767 191
rect 836 187 861 191
rect 880 187 890 191
rect 897 187 906 191
rect 959 187 996 191
rect 1015 187 1025 191
rect 1032 187 1041 191
rect -31 168 -27 187
rect -15 180 33 184
rect 43 182 47 187
rect -15 176 -11 180
rect -17 172 -11 176
rect -148 164 -103 168
rect -96 164 -27 168
rect -148 2 -144 164
rect -96 157 -92 164
rect -104 149 -100 153
rect -96 149 -92 153
rect -104 140 -100 145
rect -126 136 -111 140
rect -107 136 -100 140
rect -96 136 -89 140
rect -105 101 -98 105
rect -94 101 -87 105
rect -83 101 -60 105
rect -102 95 -98 101
rect -102 86 -98 91
rect -102 78 -98 82
rect -102 70 -98 74
rect -94 95 -90 96
rect -94 86 -90 91
rect -94 78 -90 82
rect -94 70 -90 74
rect -94 59 -90 66
rect -15 59 -11 172
rect 40 178 47 182
rect 40 170 44 178
rect 13 163 17 166
rect 13 156 17 159
rect 40 163 44 166
rect 40 156 44 159
rect 52 161 56 162
rect 13 146 17 152
rect 12 142 16 146
rect 20 142 24 146
rect 28 142 32 146
rect 36 142 40 146
rect 44 142 48 146
rect 52 142 56 157
rect 60 161 64 187
rect 130 180 173 184
rect 183 182 187 187
rect 180 178 187 182
rect 180 170 184 178
rect 60 156 64 157
rect 153 163 157 166
rect 153 156 157 159
rect 180 163 184 166
rect 180 156 184 159
rect 192 161 196 162
rect 153 146 157 152
rect 60 142 64 146
rect 68 142 95 146
rect 100 142 148 146
rect 152 142 156 146
rect 160 142 164 146
rect 168 142 172 146
rect 176 142 180 146
rect 184 142 188 146
rect 192 142 196 157
rect 200 161 204 187
rect 267 180 313 184
rect 323 182 327 187
rect 320 178 327 182
rect 320 170 324 178
rect 200 156 204 157
rect 293 163 297 166
rect 293 156 297 159
rect 320 163 324 166
rect 320 156 324 159
rect 332 161 336 162
rect 293 146 297 152
rect 200 142 204 146
rect 208 142 288 146
rect 292 142 296 146
rect 300 142 304 146
rect 308 142 312 146
rect 316 142 320 146
rect 324 142 328 146
rect 332 142 336 157
rect 340 161 344 187
rect 421 180 460 184
rect 470 182 474 187
rect 467 178 474 182
rect 467 170 471 178
rect 340 156 344 157
rect 440 163 444 166
rect 440 156 444 159
rect 467 163 471 166
rect 467 156 471 159
rect 479 161 483 162
rect 440 146 444 152
rect 340 142 344 146
rect 348 142 435 146
rect 439 142 443 146
rect 447 142 451 146
rect 455 142 459 146
rect 463 142 467 146
rect 471 142 475 146
rect 479 142 483 157
rect 487 161 491 187
rect 547 180 594 184
rect 604 182 608 187
rect 601 178 608 182
rect 601 170 605 178
rect 487 156 491 157
rect 574 163 578 166
rect 574 156 578 159
rect 601 163 605 166
rect 601 156 605 159
rect 613 161 617 162
rect 574 146 578 152
rect 487 142 491 146
rect 495 142 569 146
rect 573 142 577 146
rect 581 142 585 146
rect 589 142 593 146
rect 597 142 601 146
rect 605 142 609 146
rect 613 142 617 157
rect 621 161 625 187
rect 697 180 731 184
rect 741 182 745 187
rect 738 178 745 182
rect 738 170 742 178
rect 621 156 625 157
rect 711 163 715 166
rect 711 156 715 159
rect 738 163 742 166
rect 738 156 742 159
rect 750 161 754 162
rect 711 146 715 152
rect 621 142 625 146
rect 629 142 706 146
rect 710 142 714 146
rect 718 142 722 146
rect 726 142 730 146
rect 734 142 738 146
rect 742 142 746 146
rect 750 142 754 157
rect 758 161 762 187
rect 802 180 870 184
rect 880 182 884 187
rect 877 178 884 182
rect 877 170 881 178
rect 758 156 762 157
rect 850 163 854 166
rect 850 156 854 159
rect 877 163 881 166
rect 877 156 881 159
rect 889 161 893 162
rect 850 146 854 152
rect 758 142 762 146
rect 766 142 845 146
rect 849 142 853 146
rect 857 142 861 146
rect 865 142 869 146
rect 873 142 877 146
rect 881 142 885 146
rect 889 142 893 157
rect 897 161 901 187
rect 941 180 1005 184
rect 1015 182 1019 187
rect 1012 178 1019 182
rect 1012 170 1016 178
rect 897 156 901 157
rect 985 163 989 166
rect 985 156 989 159
rect 1012 163 1016 166
rect 1012 156 1016 159
rect 1024 161 1028 162
rect 985 146 989 152
rect 897 142 901 146
rect 905 142 980 146
rect 984 142 988 146
rect 992 142 996 146
rect 1000 142 1004 146
rect 1008 142 1012 146
rect 1016 142 1020 146
rect 1024 142 1028 157
rect 1032 161 1036 187
rect 1032 156 1036 157
rect 1032 142 1036 146
rect 1040 142 1041 146
rect -127 55 -101 59
rect -94 55 -11 59
rect 5 123 126 127
rect 131 123 417 127
rect 422 123 693 127
rect 698 123 937 127
rect -127 14 -123 55
rect -94 48 -90 55
rect -102 40 -98 44
rect -94 40 -90 44
rect -102 31 -98 36
rect -114 27 -109 31
rect -105 27 -98 31
rect -94 27 -87 31
rect 5 14 10 123
rect -127 10 10 14
rect 19 107 250 111
rect 255 107 398 111
rect 403 107 832 111
rect 837 107 955 111
rect 19 2 24 107
rect -148 -2 24 2
rect 36 91 531 95
rect 536 91 669 95
rect 674 91 815 95
rect 820 91 970 95
rect 36 -8 41 91
rect -155 -12 41 -8
<< metal2 >>
rect -56 314 80 318
rect -60 261 -56 314
rect -130 140 -126 240
rect -130 63 -126 136
rect -60 214 -56 257
rect -60 152 -56 210
rect -31 276 4 280
rect -31 238 -27 276
rect -31 191 -27 234
rect -21 260 4 264
rect -21 223 -17 260
rect 76 234 80 314
rect -21 176 -17 219
rect 108 191 112 276
rect 129 198 133 292
rect -60 105 -56 148
rect 95 63 100 142
rect 126 140 130 180
rect 250 140 254 187
rect 263 184 267 260
rect 273 198 277 292
rect 410 198 414 292
rect 398 140 402 187
rect 417 140 421 180
rect 531 140 535 194
rect 543 184 547 260
rect 554 191 558 276
rect 669 140 673 194
rect 685 191 689 276
rect 798 184 802 260
rect 693 140 697 180
rect 815 140 819 194
rect 832 140 836 187
rect 937 140 941 180
rect 955 140 959 187
rect 970 140 974 194
rect 126 127 131 140
rect 250 111 255 140
rect 398 111 403 140
rect 417 127 422 140
rect 531 95 536 140
rect 669 95 674 140
rect 693 127 698 140
rect 815 95 820 140
rect 832 111 837 140
rect 937 127 942 140
rect 955 111 960 140
rect 970 95 975 140
rect -130 59 100 63
rect -130 31 -126 59
rect -130 27 -118 31
<< ntransistor >>
rect -98 249 -96 261
rect -99 145 -97 157
rect 18 152 20 170
rect 28 152 30 170
rect 37 152 39 170
rect 57 156 59 162
rect 158 152 160 170
rect 168 152 170 170
rect 177 152 179 170
rect 197 156 199 162
rect 298 152 300 170
rect 308 152 310 170
rect 317 152 319 170
rect 337 156 339 162
rect 445 152 447 170
rect 455 152 457 170
rect 464 152 466 170
rect 484 156 486 162
rect 579 152 581 170
rect 589 152 591 170
rect 598 152 600 170
rect 618 156 620 162
rect 716 152 718 170
rect 726 152 728 170
rect 735 152 737 170
rect 755 156 757 162
rect 855 152 857 170
rect 865 152 867 170
rect 874 152 876 170
rect 894 156 896 162
rect 990 152 992 170
rect 1000 152 1002 170
rect 1009 152 1011 170
rect 1029 156 1031 162
rect -97 36 -95 48
<< ptransistor >>
rect -98 279 -96 309
rect 18 209 20 224
rect 28 209 30 224
rect 37 209 39 224
rect -99 175 -97 205
rect 57 208 59 225
rect 158 209 160 224
rect 168 209 170 224
rect 177 209 179 224
rect 197 208 199 225
rect 298 209 300 224
rect 308 209 310 224
rect 317 209 319 224
rect 337 208 339 225
rect 445 209 447 224
rect 455 209 457 224
rect 464 209 466 224
rect 484 208 486 225
rect 579 209 581 224
rect 589 209 591 224
rect 598 209 600 224
rect 618 208 620 225
rect 716 209 718 224
rect 726 209 728 224
rect 735 209 737 224
rect 755 208 757 225
rect 855 209 857 224
rect 865 209 867 224
rect 874 209 876 224
rect 894 208 896 225
rect 990 209 992 224
rect 1000 209 1002 224
rect 1009 209 1011 224
rect 1029 208 1031 225
rect -97 66 -95 96
<< polycontact >>
rect -102 268 -98 272
rect 14 194 18 198
rect -103 164 -99 168
rect 24 187 28 191
rect 33 180 37 184
rect 53 187 57 191
rect 154 194 158 198
rect 164 187 168 191
rect 173 180 177 184
rect 193 187 197 191
rect 294 194 298 198
rect 304 187 308 191
rect 313 180 317 184
rect 333 187 337 191
rect 441 194 445 198
rect 451 187 455 191
rect 460 180 464 184
rect 480 187 484 191
rect 575 194 579 198
rect 585 187 589 191
rect 594 180 598 184
rect 614 187 618 191
rect 712 194 716 198
rect 722 187 726 191
rect 731 180 735 184
rect 751 187 755 191
rect 851 194 855 198
rect 861 187 865 191
rect 870 180 874 184
rect 890 187 894 191
rect 986 194 990 198
rect 996 187 1000 191
rect 1005 180 1009 184
rect 1025 187 1029 191
rect -101 55 -97 59
<< ndcontact >>
rect -103 257 -99 261
rect -103 249 -99 253
rect -95 257 -91 261
rect -95 249 -91 253
rect 13 166 17 170
rect 13 159 17 163
rect -104 153 -100 157
rect -104 145 -100 149
rect -96 153 -92 157
rect 13 152 17 156
rect 40 166 44 170
rect 40 159 44 163
rect 153 166 157 170
rect 52 157 56 161
rect 60 157 64 161
rect 153 159 157 163
rect 40 152 44 156
rect 153 152 157 156
rect 180 166 184 170
rect 180 159 184 163
rect 293 166 297 170
rect 192 157 196 161
rect 200 157 204 161
rect 293 159 297 163
rect 180 152 184 156
rect 293 152 297 156
rect 320 166 324 170
rect 320 159 324 163
rect 440 166 444 170
rect 332 157 336 161
rect 340 157 344 161
rect 440 159 444 163
rect 320 152 324 156
rect 440 152 444 156
rect 467 166 471 170
rect 467 159 471 163
rect 574 166 578 170
rect 479 157 483 161
rect 487 157 491 161
rect 574 159 578 163
rect 467 152 471 156
rect 574 152 578 156
rect 601 166 605 170
rect 601 159 605 163
rect 711 166 715 170
rect 613 157 617 161
rect 621 157 625 161
rect 711 159 715 163
rect 601 152 605 156
rect 711 152 715 156
rect 738 166 742 170
rect 738 159 742 163
rect 850 166 854 170
rect 750 157 754 161
rect 758 157 762 161
rect 850 159 854 163
rect 738 152 742 156
rect 850 152 854 156
rect 877 166 881 170
rect 877 159 881 163
rect 985 166 989 170
rect 889 157 893 161
rect 897 157 901 161
rect 985 159 989 163
rect 877 152 881 156
rect 985 152 989 156
rect 1012 166 1016 170
rect 1012 159 1016 163
rect 1024 157 1028 161
rect 1032 157 1036 161
rect 1012 152 1016 156
rect -96 145 -92 149
rect -102 44 -98 48
rect -102 36 -98 40
rect -94 44 -90 48
rect -94 36 -90 40
<< pdcontact >>
rect -103 304 -99 308
rect -103 295 -99 299
rect -103 287 -99 291
rect -103 279 -99 283
rect -95 304 -91 308
rect -95 295 -91 299
rect -95 287 -91 291
rect -95 279 -91 283
rect 13 220 17 224
rect 13 209 17 213
rect 22 220 26 224
rect 22 209 26 213
rect 32 220 36 224
rect 32 209 36 213
rect 40 220 44 224
rect 40 209 44 213
rect 52 220 56 224
rect 52 214 56 218
rect -104 200 -100 204
rect -104 191 -100 195
rect -104 183 -100 187
rect -104 175 -100 179
rect -96 200 -92 204
rect -96 191 -92 195
rect -96 183 -92 187
rect -96 175 -92 179
rect 52 208 56 212
rect 60 220 64 224
rect 60 214 64 218
rect 60 208 64 212
rect 153 220 157 224
rect 153 209 157 213
rect 162 220 166 224
rect 162 209 166 213
rect 172 220 176 224
rect 172 209 176 213
rect 180 220 184 224
rect 180 209 184 213
rect 192 220 196 224
rect 192 214 196 218
rect 192 208 196 212
rect 200 220 204 224
rect 200 214 204 218
rect 200 208 204 212
rect 293 220 297 224
rect 293 209 297 213
rect 302 220 306 224
rect 302 209 306 213
rect 312 220 316 224
rect 312 209 316 213
rect 320 220 324 224
rect 320 209 324 213
rect 332 220 336 224
rect 332 214 336 218
rect 332 208 336 212
rect 340 220 344 224
rect 340 214 344 218
rect 340 208 344 212
rect 440 220 444 224
rect 440 209 444 213
rect 449 220 453 224
rect 449 209 453 213
rect 459 220 463 224
rect 459 209 463 213
rect 467 220 471 224
rect 467 209 471 213
rect 479 220 483 224
rect 479 214 483 218
rect 479 208 483 212
rect 487 220 491 224
rect 487 214 491 218
rect 487 208 491 212
rect 574 220 578 224
rect 574 209 578 213
rect 583 220 587 224
rect 583 209 587 213
rect 593 220 597 224
rect 593 209 597 213
rect 601 220 605 224
rect 601 209 605 213
rect 613 220 617 224
rect 613 214 617 218
rect 613 208 617 212
rect 621 220 625 224
rect 621 214 625 218
rect 621 208 625 212
rect 711 220 715 224
rect 711 209 715 213
rect 720 220 724 224
rect 720 209 724 213
rect 730 220 734 224
rect 730 209 734 213
rect 738 220 742 224
rect 738 209 742 213
rect 750 220 754 224
rect 750 214 754 218
rect 750 208 754 212
rect 758 220 762 224
rect 758 214 762 218
rect 758 208 762 212
rect 850 220 854 224
rect 850 209 854 213
rect 859 220 863 224
rect 859 209 863 213
rect 869 220 873 224
rect 869 209 873 213
rect 877 220 881 224
rect 877 209 881 213
rect 889 220 893 224
rect 889 214 893 218
rect 889 208 893 212
rect 897 220 901 224
rect 897 214 901 218
rect 897 208 901 212
rect 985 220 989 224
rect 985 209 989 213
rect 994 220 998 224
rect 994 209 998 213
rect 1004 220 1008 224
rect 1004 209 1008 213
rect 1012 220 1016 224
rect 1012 209 1016 213
rect 1024 220 1028 224
rect 1024 214 1028 218
rect 1024 208 1028 212
rect 1032 220 1036 224
rect 1032 214 1036 218
rect 1032 208 1036 212
rect -102 91 -98 95
rect -102 82 -98 86
rect -102 74 -98 78
rect -102 66 -98 70
rect -94 91 -90 95
rect -94 82 -90 86
rect -94 74 -90 78
rect -94 66 -90 70
<< m2contact >>
rect -60 314 -56 318
rect 129 292 133 296
rect 273 292 277 296
rect 410 292 414 296
rect -60 257 -56 261
rect -130 240 -126 244
rect -31 234 -27 238
rect -21 219 -17 223
rect -60 210 -56 214
rect 4 276 8 280
rect 108 276 112 280
rect 554 276 558 280
rect 685 276 689 280
rect 4 260 8 264
rect 263 260 267 264
rect 543 260 547 264
rect 798 260 802 264
rect 76 230 80 234
rect 129 194 133 198
rect 273 194 277 198
rect 410 194 414 198
rect 531 194 535 198
rect 669 194 673 198
rect 815 194 819 198
rect 970 194 974 198
rect -31 187 -27 191
rect 108 187 112 191
rect 250 187 254 191
rect 398 187 402 191
rect 554 187 558 191
rect 685 187 689 191
rect 832 187 836 191
rect 955 187 959 191
rect -21 172 -17 176
rect -60 148 -56 152
rect -130 136 -126 140
rect -60 101 -56 105
rect 126 180 130 184
rect 95 142 100 146
rect 263 180 267 184
rect 417 180 421 184
rect 543 180 547 184
rect 693 180 697 184
rect 798 180 802 184
rect 937 180 941 184
rect 126 123 131 127
rect 417 123 422 127
rect 693 123 698 127
rect 937 123 942 127
rect -118 27 -114 31
rect 250 107 255 111
rect 398 107 403 111
rect 832 107 837 111
rect 955 107 960 111
rect 531 91 536 95
rect 669 91 674 95
rect 815 91 820 95
rect 970 91 975 95
<< psubstratepcontact >>
rect -110 240 -106 244
rect -99 240 -95 244
rect -88 240 -84 244
rect 8 142 12 146
rect 16 142 20 146
rect 24 142 28 146
rect 32 142 36 146
rect 40 142 44 146
rect 48 142 52 146
rect 56 142 60 146
rect 64 142 68 146
rect 148 142 152 146
rect 156 142 160 146
rect 164 142 168 146
rect 172 142 176 146
rect 180 142 184 146
rect 188 142 192 146
rect 196 142 200 146
rect 204 142 208 146
rect 288 142 292 146
rect 296 142 300 146
rect 304 142 308 146
rect 312 142 316 146
rect 320 142 324 146
rect 328 142 332 146
rect 336 142 340 146
rect 344 142 348 146
rect 435 142 439 146
rect 443 142 447 146
rect 451 142 455 146
rect 459 142 463 146
rect 467 142 471 146
rect 475 142 479 146
rect 483 142 487 146
rect 491 142 495 146
rect 569 142 573 146
rect 577 142 581 146
rect 585 142 589 146
rect 593 142 597 146
rect 601 142 605 146
rect 609 142 613 146
rect 617 142 621 146
rect 625 142 629 146
rect 706 142 710 146
rect 714 142 718 146
rect 722 142 726 146
rect 730 142 734 146
rect 738 142 742 146
rect 746 142 750 146
rect 754 142 758 146
rect 762 142 766 146
rect 845 142 849 146
rect 853 142 857 146
rect 861 142 865 146
rect 869 142 873 146
rect 877 142 881 146
rect 885 142 889 146
rect 893 142 897 146
rect 901 142 905 146
rect 980 142 984 146
rect 988 142 992 146
rect 996 142 1000 146
rect 1004 142 1008 146
rect 1012 142 1016 146
rect 1020 142 1024 146
rect 1028 142 1032 146
rect 1036 142 1040 146
rect -111 136 -107 140
rect -100 136 -96 140
rect -89 136 -85 140
rect -109 27 -105 31
rect -98 27 -94 31
rect -87 27 -83 31
<< nsubstratencontact >>
rect -110 314 -106 318
rect -99 314 -95 318
rect -88 314 -84 318
rect 8 230 12 234
rect 16 230 20 234
rect 24 230 28 234
rect 32 230 36 234
rect 40 230 44 234
rect 48 230 52 234
rect 56 230 60 234
rect 64 230 68 234
rect 148 230 152 234
rect 156 230 160 234
rect 164 230 168 234
rect 172 230 176 234
rect 180 230 184 234
rect 188 230 192 234
rect 196 230 200 234
rect 204 230 208 234
rect 288 230 292 234
rect 296 230 300 234
rect 304 230 308 234
rect 312 230 316 234
rect 320 230 324 234
rect 328 230 332 234
rect 336 230 340 234
rect 344 230 348 234
rect 435 230 439 234
rect 443 230 447 234
rect 451 230 455 234
rect 459 230 463 234
rect 467 230 471 234
rect 475 230 479 234
rect 483 230 487 234
rect 491 230 495 234
rect 569 230 573 234
rect 577 230 581 234
rect 585 230 589 234
rect 593 230 597 234
rect 601 230 605 234
rect 609 230 613 234
rect 617 230 621 234
rect 625 230 629 234
rect 706 230 710 234
rect 714 230 718 234
rect 722 230 726 234
rect 730 230 734 234
rect 738 230 742 234
rect 746 230 750 234
rect 754 230 758 234
rect 762 230 766 234
rect 845 230 849 234
rect 853 230 857 234
rect 861 230 865 234
rect 869 230 873 234
rect 877 230 881 234
rect 885 230 889 234
rect 893 230 897 234
rect 901 230 905 234
rect 980 230 984 234
rect 988 230 992 234
rect 996 230 1000 234
rect 1004 230 1008 234
rect 1012 230 1016 234
rect 1020 230 1024 234
rect 1028 230 1032 234
rect 1036 230 1040 234
rect -111 210 -107 214
rect -100 210 -96 214
rect -89 210 -85 214
rect -109 101 -105 105
rect -98 101 -94 105
rect -87 101 -83 105
<< labels >>
rlabel metal1 69 187 69 191 1 out0
rlabel metal1 209 187 209 191 1 out1
rlabel metal1 349 187 349 191 1 out2
rlabel metal1 496 187 496 191 1 out3
rlabel metal1 630 187 630 191 1 out4
rlabel metal1 767 187 767 191 1 out5
rlabel metal1 906 187 906 191 1 out6
rlabel metal1 1041 187 1041 191 1 out7
rlabel metal1 1041 230 1041 234 1 vdd
rlabel metal1 1041 142 1041 146 1 gnd
rlabel metal1 -118 268 -118 272 1 a
rlabel metal1 -116 164 -116 168 1 b
rlabel metal1 -114 55 -114 59 1 c
rlabel metal1 -71 55 -71 59 1 c_out
rlabel metal1 -77 164 -77 168 1 b_out
rlabel metal1 -78 268 -78 272 1 a_out
<< end >>
